   
    parameter PROC_NUM = 47;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    reg stop_report_path;
    reg [PROC_NUM - 1:0] reported_proc;
    integer i;
    integer fp;

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            reported_proc <= 'b0;
        end
        else if (CS_fsm == ST_DL_REPORT) begin
            reported_proc <= reported_proc | dl_in_vec;
        end
        else if (CS_fsm == ST_DL_DETECTED) begin
            reported_proc <= 'b0;
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            stop_report_path <= 1'b0;
        end
        else if (CS_fsm == ST_DL_REPORT && (|(dl_in_vec & reported_proc))) begin
            stop_report_path <= 1'b1;
        end
        else if (CS_fsm == ST_IDLE) begin
            stop_report_path <= 1'b0;
        end
    end

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end

    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if ((dl_detect_reg != dl_done_reg) && stop_report_path == 1'b0) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                // avoid report deadlock ring.
                else if (|(dl_in_vec & reported_proc)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && ((dl_detect_reg == dl_done_reg) || (stop_report_path == 1'b1))) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [1592:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0";
                end
                1 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0";
                end
                2 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0";
                end
                3 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0";
                end
                4 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0";
                end
                5 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0";
                end
                6 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0";
                end
                7 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0";
                end
                8 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0";
                end
                9 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0";
                end
                10 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0";
                end
                11 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0";
                end
                12 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0";
                end
                13 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0";
                end
                14 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0";
                end
                15 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0";
                end
                16 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0";
                end
                17 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0";
                end
                18 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0";
                end
                19 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0";
                end
                20 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0";
                end
                21 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0";
                end
                22 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0";
                end
                23 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0";
                end
                24 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0";
                end
                25 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0";
                end
                26 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0";
                end
                27 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0";
                end
                28 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0";
                end
                29 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0";
                end
                30 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0";
                end
                31 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0";
                end
                32 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0";
                end
                33 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0";
                end
                34 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0";
                end
                35 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0";
                end
                36 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0";
                end
                37 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0";
                end
                38 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0";
                end
                39 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0";
                end
                40 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0";
                end
                41 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0";
                end
                42 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0";
                end
                43 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0";
                end
                44 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0";
                end
                45 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0";
                end
                46 : begin
                    proc_path = "Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [1592:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [1592:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [1656:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'
                    case(index2)
                    2: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Block_entry_split_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready} input_sync}
                        if ((ap_sync_Block_entry_split_proc_U0_ap_ready & Block_entry_split_proc_U0.ap_idle & ~ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'");
                        end
                    end
                    18: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Block_entry_split_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready} input_sync}
                        if ((ap_sync_Block_entry_split_proc_U0_ap_ready & Block_entry_split_proc_U0.ap_idle & ~ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'");
                        end
                    end
                    endcase
                end
                1 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
                    case(index2)
                    0: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_out_tmp_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_out_tmp_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Process_N_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_out_tmp_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_out_tmp_channel_U.if_empty_n & Process_N_U0.ap_idle & ~nCols_assign_out_tmp_channel_U.if_write)) begin
                            if (~nCols_assign_out_tmp_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_out_tmp_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_out_tmp_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_out_tmp_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_out_tmp_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_out_tmp_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_out_tmp_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_out_tmp_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Process_N_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_out_tmp_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_out_tmp_channel_U.if_empty_n & Process_N_U0.ap_idle & ~nRows_assign_out_tmp_channel_U.if_write)) begin
                            if (~nRows_assign_out_tmp_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_out_tmp_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_out_tmp_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_out_tmp_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_out_tmp_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_out_tmp_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                2 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'
                    case(index2)
                    46: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.dPrimalInfeasRes_blk_n data_FIFO} {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_noScaled_fu_72.twoNorm_U0.dPrimalInfeasRes_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.dPrimalInfeasRes_blk_n) | (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_noScaled_fu_72.twoNorm_U0.dPrimalInfeasRes_blk_n)) begin
                            if (~dPrimalInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dPrimalInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.real_start & (trans_in_cnt_13 == trans_out_cnt_13) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_read} start_FIFO}
                        if ((~start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.real_start & (trans_in_cnt_13 == trans_out_cnt_13) & ~start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0',");
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c2_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c2_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c2_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~nRows_assign_c2_channel_U.if_write)) begin
                            if (~nRows_assign_c2_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c2_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c3_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~nCols_assign_c3_channel_U.if_write)) begin
                            if (~nCols_assign_c3_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c3_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Block_entry_split_proc_U0_ap_ready} input_sync}
                        if ((ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~ap_sync_Block_entry_split_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                        end
                    end
                    18: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready} input_sync}
                        if ((ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.ap_idle & ~ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'");
                        end
                    end
                    endcase
                end
                3 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
                    case(index2)
                    11: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0',");
                        end
                    end
                    10: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c5_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c5_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0',");
                        end
                    end
                    9: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c6_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c6_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0',");
                        end
                    end
                    8: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c7_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.inverse_dScale_c7_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0',");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                4 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
                    case(index2)
                    8: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.grp_loadDDR_data_Pipeline_loadDDR_data_fu_84.dualInfeasRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.grp_loadDDR_data_Pipeline_loadDDR_data_fu_84.dualInfeasRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.nRows_assign_c1_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.nRows_assign_c1_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c2_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c2_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c2_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~nRows_assign_c2_channel_U.if_write)) begin
                            if (~nRows_assign_c2_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c2_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c2_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                5 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
                    case(index2)
                    9: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.grp_loadDDR_data_15_Pipeline_loadDDR_data_fu_84.dualInfeasLbRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.grp_loadDDR_data_15_Pipeline_loadDDR_data_fu_84.dualInfeasLbRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.nCols_assign_c4_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.nCols_assign_c4_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c3_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~nCols_assign_c3_channel_U.if_write)) begin
                            if (~nCols_assign_c3_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c3_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                6 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
                    case(index2)
                    10: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.grp_loadDDR_data_16_Pipeline_loadDDR_data_fu_84.dualInfeasUbRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.grp_loadDDR_data_16_Pipeline_loadDDR_data_fu_84.dualInfeasUbRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.nCols_assign_c3_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.nCols_assign_c3_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c3_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~nCols_assign_c3_channel_U.if_write)) begin
                            if (~nCols_assign_c3_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c3_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                7 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
                    case(index2)
                    11: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.grp_loadDDR_data_17_Pipeline_loadDDR_data_fu_84.dualInfeasConstr_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.grp_loadDDR_data_17_Pipeline_loadDDR_data_fu_84.dualInfeasConstr_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.nCols_assign_c2_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.nCols_assign_c2_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c3_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~nCols_assign_c3_channel_U.if_write)) begin
                            if (~nCols_assign_c3_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c3_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                8 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'
                    case(index2)
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.inverse_dScale_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.inverse_dScale_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_12_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0',");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.grp_scaleVector_12_Pipeline_scale_vector_fu_60.dualInfeasRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.grp_scaleVector_12_Pipeline_scale_vector_fu_60.dualInfeasRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.nRows_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.nRows_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.grp_scaleVector_12_Pipeline_scale_vector_fu_60.dualInfeasRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.grp_scaleVector_12_Pipeline_scale_vector_fu_60.dualInfeasRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.nRows_assign_c_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.nRows_assign_c_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0',");
                        end
                    end
                    endcase
                end
                9 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'
                    case(index2)
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.inverse_dScale_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.inverse_dScale_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_13_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0',");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.grp_scaleVector_13_Pipeline_scale_vector_fu_48.dualInfeasLbRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.grp_scaleVector_13_Pipeline_scale_vector_fu_48.dualInfeasLbRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.grp_scaleVector_13_Pipeline_scale_vector_fu_48.dualInfeasLbRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.grp_scaleVector_13_Pipeline_scale_vector_fu_48.dualInfeasLbRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0',");
                        end
                    end
                    endcase
                end
                10 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'
                    case(index2)
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.inverse_dScale_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.inverse_dScale_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_14_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0',");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.grp_scaleVector_14_Pipeline_scale_vector_fu_48.dualInfeasUbRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.grp_scaleVector_14_Pipeline_scale_vector_fu_48.dualInfeasUbRay_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.grp_scaleVector_14_Pipeline_scale_vector_fu_48.dualInfeasUbRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0.grp_scaleVector_14_Pipeline_scale_vector_fu_48.dualInfeasUbRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'
                    case(index2)
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.inverse_dScale_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.inverse_dScale_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.inverse_dScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_scaleVector_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0',");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.grp_scaleVector_Pipeline_scale_vector_fu_60.dualInfeasConstr_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.grp_scaleVector_Pipeline_scale_vector_fu_60.dualInfeasConstr_fifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.grp_scaleVector_Pipeline_scale_vector_fu_60.dualInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.grp_scaleVector_Pipeline_scale_vector_fu_60.dualInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.nCols_assign_c_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0.nCols_assign_c_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                12 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'
                    case(index2)
                    8: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.consumer_U0.grp_consumer_Pipeline_VITIS_LOOP_15_1_fu_36.dualInfeasRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.consumer_U0.grp_consumer_Pipeline_VITIS_LOOP_15_1_fu_36.dualInfeasRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.consumer_U0.nRows_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.consumer_U0.nRows_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_consumer_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_12_U0',");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_20 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_done} output_sync}
                        if ((ap_done_reg_20 & Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_done & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                        end
                    end
                    endcase
                end
                13 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'
                    case(index2)
                    11: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasLbRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasLbRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasLbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.start_for_axpy_2fused_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_13_U0',");
                        end
                    end
                    10: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasUbRay_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasUbRay_SVfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scaleVector_14_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasUbRay_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasConstr_axpyfifo_i_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0.grp_axpy_2fused_Pipeline_axpy_2fused_fu_42.dualInfeasConstr_axpyfifo_i_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                14 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
                    case(index2)
                    13: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.dualInfeasConstr_axpyfifo_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.dualInfeasConstr_axpyfifo_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.axpy_2fused_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.dualInfeasConstr_axpyfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.dPrimalInfeasRes_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.dPrimalInfeasRes_blk_n)) begin
                            if (~dPrimalInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dPrimalInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c3_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c3_channel_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~nCols_assign_c3_channel_U.if_write)) begin
                            if (~nCols_assign_c3_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c3_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c3_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_entry_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.entry_proc_U0'");
                        end
                    end
                    4: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_U0'");
                        end
                    end
                    5: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_15_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_15_U0'");
                        end
                    end
                    6: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_16_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_16_U0'");
                        end
                    end
                    7: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready} input_sync}
                        if ((Compute_Primal_Infeasibility_stage2_U0.ap_sync_scale_and_twoNorm_U0_ap_ready & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.ap_sync_loadDDR_data_17_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.loadDDR_data_17_U0'");
                        end
                    end
                    12: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_6 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_done} output_sync}
                        if ((ap_done_reg_6 & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.ap_done & ~Compute_Primal_Infeasibility_stage2_U0.consumer_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.consumer_U0'");
                        end
                    end
                    endcase
                end
                15 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'
                    case(index2)
                    16: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.grp_loadDDR_data_22_Pipeline_loadDDR_data_fu_84.colScale_fifo_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.grp_loadDDR_data_22_Pipeline_loadDDR_data_fu_84.colScale_fifo_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.n_c1_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.n_c1_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0',");
                        end
                    end
                    endcase
                end
                16 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'
                    case(index2)
                    15: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.colScale_fifo_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.colScale_fifo_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.colScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.n_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.n_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_edot_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.loadDDR_data_22_U0',");
                        end
                    end
                    17: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.temp_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.grp_edot_Pipeline_edot_fu_52.temp_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.n_c_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.n_c_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_read} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_full_n & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.ap_start & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0',");
                        end
                    end
                    endcase
                end
                17 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0'
                    case(index2)
                    16: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.grp_twoNorm_23_Pipeline_twoNorm_fu_55.temp_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.grp_twoNorm_23_Pipeline_twoNorm_fu_55.temp_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.n_blk_n data_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.n_blk_n)) begin
                            if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_write} start_FIFO}
                        if ((~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_empty_n & Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.twoNorm_23_U0.ap_idle & ~Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.start_for_twoNorm_23_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0.grp_scale_and_twoNorm_Scaled_fu_58.edot_U0',");
                        end
                    end
                    endcase
                end
                18 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'
                    case(index2)
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~nRows_assign_c_channel_U.if_write)) begin
                            if (~nRows_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.dDualInfeasRes_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.dDualInfeasRes_blk_n)) begin
                            if (~dDualInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dDualInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    0: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Block_entry_split_proc_U0_ap_ready} input_sync}
                        if ((ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~ap_sync_Block_entry_split_proc_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_proc_U0'");
                        end
                    end
                    2: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready} input_sync}
                        if ((ap_sync_Compute_Dual_Infeasibility_stage2_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.ap_idle & ~ap_sync_Compute_Primal_Infeasibility_stage2_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'");
                        end
                    end
                    endcase
                end
                19 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
                    case(index2)
                    23: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.inverse_pScale_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.inverse_pScale_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0',");
                        end
                    end
                    22: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.inverse_pScale_c1_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.inverse_pScale_c1_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0',");
                        end
                    end
                    20: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                        end
                    end
                    21: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                        end
                    end
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                        end
                    end
                    endcase
                end
                20 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
                    case(index2)
                    22: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.grp_loadDDR_data_18_Pipeline_loadDDR_data_fu_84.primalInfeasRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.grp_loadDDR_data_18_Pipeline_loadDDR_data_fu_84.primalInfeasRay_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.nCols_assign_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.nCols_assign_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                        end
                    end
                    21: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                        end
                    end
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                        end
                    end
                    endcase
                end
                21 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
                    case(index2)
                    23: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.grp_loadDDR_data_19_Pipeline_loadDDR_data_fu_84.primalINfeasConstr_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.grp_loadDDR_data_19_Pipeline_loadDDR_data_fu_84.primalINfeasConstr_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.nRows_assign_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.nRows_assign_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~nRows_assign_c_channel_U.if_write)) begin
                            if (~nRows_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                        end
                    end
                    20: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                        end
                    end
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                        end
                    end
                    endcase
                end
                22 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
                    case(index2)
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.inverse_pScale_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.inverse_pScale_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_2out_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0',");
                        end
                    end
                    20: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0.grp_scaleVector_2out_Pipeline_scale_vector_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                23 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'
                    case(index2)
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.inverse_pScale_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.inverse_pScale_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.inverse_pScale_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.start_for_scaleVector_1_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0',");
                        end
                    end
                    21: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalINfeasConstr_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalINfeasConstr_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalINfeasConstr_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.nRows_assign_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.nRows_assign_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.nRows_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0.grp_scaleVector_1_Pipeline_scale_vector_fu_48.primalInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                24 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
                    case(index2)
                    23: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~nRows_assign_c_channel_U.if_write)) begin
                            if (~nRows_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_done & ap_done_reg_10 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_done & ap_done_reg_10 & ~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                        end
                    end
                    20: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                        end
                    end
                    21: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                        end
                    end
                    endcase
                end
                25 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'
                    case(index2)
                    23: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasConstr_SVfifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasConstr_SVfifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasConstr_SVfifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasBound_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.primalInfeasBound_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_projNeg28_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_scale_and_twoNormSquared29_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_projNeg28_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_scale_and_twoNormSquared29_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'");
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0.ap_idle & ~nRows_assign_c_channel_U.if_write)) begin
                            if (~nRows_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                26 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'
                    case(index2)
                    25: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_noScaled_fu_72.twoNormSquared_10_U0.grp_twoNormSquared_10_Pipeline_accum_loop_fu_153.primalInfeasBound_fifo_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_noScaled_fu_72.twoNormSquared_10_U0.grp_twoNormSquared_10_Pipeline_accum_loop_fu_153.primalInfeasBound_fifo_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.primalInfeasBound_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_scale_and_twoNormSquared29_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_projNeg28_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_scale_and_twoNormSquared29_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.ap_sync_projNeg28_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.projNeg28_U0'");
                        end
                    end
                    45: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_done & ap_done_reg_12 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_done & ap_done_reg_12 & ~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nRows_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nRows_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.ap_idle & ~nRows_assign_c_channel_U.if_write)) begin
                            if (~nRows_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nRows_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nRows_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                27 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'
                    case(index2)
                    28: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.grp_loadDDR_data_24_Pipeline_loadDDR_data_fu_84.rowScale_fifo_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.grp_loadDDR_data_24_Pipeline_loadDDR_data_fu_84.rowScale_fifo_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.n_c1_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.n_c1_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.real_start & (trans_in_cnt_6 == trans_out_cnt_6) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0.real_start & (trans_in_cnt_6 == trans_out_cnt_6) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0',");
                        end
                    end
                    endcase
                end
                28 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'
                    case(index2)
                    27: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.grp_edot_11_Pipeline_edot_fu_52.rowScale_fifo_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.grp_edot_11_Pipeline_edot_fu_52.rowScale_fifo_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.rowScale_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_edot_11_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.loadDDR_data_24_U0',");
                        end
                    end
                    29: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.grp_edot_11_Pipeline_edot_fu_52.temp_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.grp_edot_11_Pipeline_edot_fu_52.temp_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.n_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.n_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.real_start & (trans_in_cnt_7 == trans_out_cnt_7) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0.real_start & (trans_in_cnt_7 == trans_out_cnt_7) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0',");
                        end
                    end
                    endcase
                end
                29 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0'
                    case(index2)
                    28: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.grp_twoNormSquared_Pipeline_accum_loop_fu_163.temp_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.grp_twoNormSquared_Pipeline_accum_loop_fu_163.temp_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.temp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.n_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.twoNormSquared_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.start_for_twoNormSquared_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0.grp_scale_and_twoNormSquared_Scaled_fu_58.edot_11_U0',");
                        end
                    end
                    endcase
                end
                30 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
                    case(index2)
                    22: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_done & ap_done_reg_13 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_done & ap_done_reg_13 & ~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_done & ap_done_reg_13 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_done & ap_done_reg_13 & ~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_entry_proc31_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.entry_proc31_U0'");
                        end
                    end
                    20: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_18_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_18_U0'");
                        end
                    end
                    21: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_loadDDR_data_19_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.loadDDR_data_19_U0'");
                        end
                    end
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Bound_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.ap_sync_Primal_Constr_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                        end
                    end
                    endcase
                end
                31 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
                    case(index2)
                    22: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasRay_SVfifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasBound_fifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.grp_projNeg_221_Pipeline_projNeg_fu_50.primalInfeasBound_fifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.nCols_assign_c1_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.nCols_assign_c1_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0',");
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                        end
                    end
                    33: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                        end
                    end
                    34: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                        end
                    end
                    endcase
                end
                32 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
                    case(index2)
                    22: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasRay_SVfifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.scaleVector_2out_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.primalInfeasRay_SVfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasBound_fifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.grp_projPos22_Pipeline_projPos_fu_50.primalInfeasBound_fifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.nCols_assign_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.nCols_assign_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0',");
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                        end
                    end
                    33: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                        end
                    end
                    34: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                        end
                    end
                    endcase
                end
                33 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
                    case(index2)
                    35: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.hasLower_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.hasLower_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                        end
                    end
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                        end
                    end
                    34: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                        end
                    end
                    endcase
                end
                34 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
                    case(index2)
                    36: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.hasUpper_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.hasUpper_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                        end
                    end
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                        end
                    end
                    33: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                        end
                    end
                    endcase
                end
                35 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'
                    case(index2)
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.primalInfeasBound_fifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.primalInfeasBound_fifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_325_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0',");
                        end
                    end
                    33: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.hasLower_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.hasLower_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasLower_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.primalInfeasBound_edotfifo_lb_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0.grp_edot_325_Pipeline_edot_fu_40.primalInfeasBound_edotfifo_lb_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                36 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'
                    case(index2)
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.primalInfeasBound_fifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.primalInfeasBound_fifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_fifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.nCols_assign_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.nCols_assign_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.nCols_assign_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.start_for_edot_426_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0',");
                        end
                    end
                    34: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.hasUpper_fifo_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.hasUpper_fifo_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.hasUpper_fifo_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.primalInfeasBound_edotfifo_ub_i_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0.grp_edot_426_Pipeline_edot_fu_40.primalInfeasBound_edotfifo_ub_i_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                37 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
                    case(index2)
                    35: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.primalInfeasBound_edotfifo_lb_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.primalInfeasBound_edotfifo_lb_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_325_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_lb_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.primalInfeasBound_edotfifo_ub_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.primalInfeasBound_edotfifo_ub_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.edot_426_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.primalInfeasBound_edotfifo_ub_i_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_done & ap_done_reg_18 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_done & ap_done_reg_18 & ~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_done & ap_done_reg_18 & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_read} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_done & ap_done_reg_18 & ~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_read)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.nCols_assign_c_channel_U.if_write} TLF_FIFO}
                        if ((~nCols_assign_c_channel_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~nCols_assign_c_channel_U.if_write)) begin
                            if (~nCols_assign_c_channel_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~nCols_assign_c_channel_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Process_N_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.nCols_assign_c_channel_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projNeg_221_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projNeg_221_U0'");
                        end
                    end
                    32: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_projPos22_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.projPos22_U0'");
                        end
                    end
                    33: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2023_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2023_U0'");
                        end
                    end
                    34: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready} input_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_scale_and_twoNormSquared_for_lub27_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.ap_sync_loadDDR_data_2124_U0_ap_ready)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.loadDDR_data_2124_U0'");
                        end
                    end
                    endcase
                end
                38 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'
                    case(index2)
                    39: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.grp_loadDDR_data_special_Pipeline_loadDDR_data_fu_96.colScale_fifo_lb_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.grp_loadDDR_data_special_Pipeline_loadDDR_data_fu_96.colScale_fifo_lb_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.nCols_c3_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.nCols_c3_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.real_start & (trans_in_cnt_10 == trans_out_cnt_10) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.real_start & (trans_in_cnt_10 == trans_out_cnt_10) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0',");
                        end
                    end
                    40: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.grp_loadDDR_data_special_Pipeline_loadDDR_data_fu_96.colScale_fifo_ub_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.grp_loadDDR_data_special_Pipeline_loadDDR_data_fu_96.colScale_fifo_ub_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.nCols_c2_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.nCols_c2_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.real_start & (trans_in_cnt_10 == trans_out_cnt_10) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0.real_start & (trans_in_cnt_10 == trans_out_cnt_10) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0',");
                        end
                    end
                    endcase
                end
                39 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'
                    case(index2)
                    38: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.colScale_fifo_lb_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.colScale_fifo_lb_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_7_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0',");
                        end
                    end
                    41: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.temp_lb_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.grp_ediv_7_Pipeline_ediv_fu_52.temp_lb_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.nCols_c1_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.nCols_c1_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.real_start & (trans_in_cnt_11 == trans_out_cnt_11) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0.real_start & (trans_in_cnt_11 == trans_out_cnt_11) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0',");
                        end
                    end
                    endcase
                end
                40 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'
                    case(index2)
                    38: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.colScale_fifo_ub_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.colScale_fifo_ub_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.colScale_fifo_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_ediv_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.loadDDR_data_special_U0',");
                        end
                    end
                    42: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.temp_ub_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.grp_ediv_Pipeline_ediv_fu_52.temp_ub_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.nCols_c_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.nCols_c_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_full_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.ap_start & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.real_start & (trans_in_cnt_12 == trans_out_cnt_12) & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_read} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_full_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.ap_start & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0.real_start & (trans_in_cnt_12 == trans_out_cnt_12) & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_read)) begin
                            $display("//      Blocked by full output start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0',");
                        end
                    end
                    endcase
                end
                41 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'
                    case(index2)
                    39: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.grp_twoNormSquared_8_Pipeline_accum_loop_fu_163.temp_lb_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.grp_twoNormSquared_8_Pipeline_accum_loop_fu_163.temp_lb_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_lb_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_8_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_7_U0',");
                        end
                    end
                    42: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_21 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_done} output_sync}
                        if ((ap_done_reg_21 & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_done & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'");
                        end
                    end
                    endcase
                end
                42 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0'
                    case(index2)
                    40: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.grp_twoNormSquared_9_Pipeline_accum_loop_fu_163.temp_ub_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.grp_twoNormSquared_9_Pipeline_accum_loop_fu_163.temp_ub_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.temp_ub_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.n_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.n_blk_n)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.nCols_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_write} start_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.start_for_twoNormSquared_9_U0_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.ediv_U0',");
                        end
                    end
                    41: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'
// for dep channel '' info is :
// blk sig is {{ap_done_reg_22 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_done} output_sync}
                        if ((ap_done_reg_22 & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_9_U0.ap_done & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0.ap_done)) begin
                            $display("//      Blocked by output sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_Scaled_fu_62.twoNormSquared_8_U0'");
                        end
                    end
                    endcase
                end
                43 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0'
                    case(index2)
                    44: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_5_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_6_U0_ap_ready} input_sync} {{ap_done_reg_23 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_done} output_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_5_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_6_U0_ap_ready) | (ap_done_reg_23 & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_done & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_done)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0'");
                        end
                    end
                    endcase
                end
                44 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0'
                    case(index2)
                    43: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0'
// for dep channel '' info is :
// blk sig is {{Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_6_U0_ap_ready & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_5_U0_ap_ready} input_sync} {{ap_done_reg_24 & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_done & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_done} output_sync}
                        if ((Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_6_U0_ap_ready & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.ap_sync_twoNormSquared_5_U0_ap_ready) | (ap_done_reg_24 & Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_6_U0.ap_done & ~Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0.ap_done)) begin
                            $display("//      Blocked by input sync logic with process : 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0.grp_scale_and_twoNormSquared_for_lub_noScaled_fu_80.twoNormSquared_5_U0'");
                        end
                    end
                    endcase
                end
                45 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
                    case(index2)
                    24: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Constr_U0.scale_and_twoNormSquared29_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pConstrResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundUbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_write} TLF_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n & Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.ap_idle & ~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_write)) begin
                            if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.Primal_Bound_U0.scale_and_twoNormSquared_for_lub27_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.pBoundLbResSq_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.dDualInfeasRes_blk_n data_FIFO}
                        if ((~Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0.dDualInfeasRes_blk_n)) begin
                            if (~dDualInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dDualInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                46 : begin // for proc 'Infeasi_Res_S2_Infeasi_Res_S2.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0'
                    case(index2)
                    2: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dPrimalInfeasRes_blk_n data_FIFO}
                        if ((~Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dPrimalInfeasRes_blk_n)) begin
                            if (~dPrimalInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dPrimalInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U' info is :
// blk sig is {{~Infeasi_Res_S2_Infeasi_Res_S2_inst.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_empty_n & Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.ap_idle & ~Infeasi_Res_S2_Infeasi_Res_S2_inst.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_write} start_FIFO}
                        if ((~start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_empty_n & Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.ap_idle & ~start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U.if_write)) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.start_for_Block_entry_split_split_split_split_split_split_split_split_split_pbkb_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0',");
                        end
                    end
                    14: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dPrimalInfeasRes_blk_n data_FIFO}
                        if ((~Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dPrimalInfeasRes_blk_n)) begin
                            if (~dPrimalInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dPrimalInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Primal_Infeasibility_stage2_U0.scale_and_twoNorm_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dPrimalInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dDualInfeasRes_blk_n data_FIFO}
                        if ((~Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dDualInfeasRes_blk_n)) begin
                            if (~dDualInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dDualInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin //  for dep proc 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'
// for dep channel 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' info is :
// blk sig is {~Infeasi_Res_S2_Infeasi_Res_S2_inst.Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dDualInfeasRes_blk_n data_FIFO}
                        if ((~Block_entry_split_split_split_split_split_split_split_split_split_proc1_U0.dDualInfeasRes_blk_n)) begin
                            if (~dDualInfeasRes_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' written by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~dDualInfeasRes_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U' read by process 'Infeasi_Res_S2_Infeasi_Res_S2.Compute_Dual_Infeasibility_stage2_U0.add3_Sqrt_U0'");
                                $fdisplay(fp, "Dependence_Channel_path Infeasi_Res_S2_Infeasi_Res_S2.dDualInfeasRes_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg && stop_report_path == 1'b0) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg)) & ~(|(reported_proc & dl_in_vec))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else if (~(|(dl_in_vec)))begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
